typedef uvm_sequencer #(encoder_transaction) encoder_sequencer;