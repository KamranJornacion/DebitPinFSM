interface encoder_if;
  logic [3:0] in;
  logic[1:0] out;
   
endinterface